`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    07:34:31 06/08/2025 
// Design Name: 
// Module Name:    FormatTiming 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module FormatTiming(
	input [2:0] GMode,
	input FrameFormat,
	input AnG,
	input Clk,
	output PixelClk,
	output reg HSn,
	output reg FSn,
	output BackPorch,
	output active,
	output Load,
	output [3:0] alphaRow,
	output DA0
   );

	wire activeRow;
	wire [9:0] frameTopRow;
	wire [9:0] frameBottomRow;
	wire [9:0] frameAllRows;
	wire slowMode;
	reg u_da0;
	reg hBlank;
	reg vBlank;

// horizontal beam counter using gclk for frame timing accuracy
	wire colReset;
	reg [8:0] colCounter;
	// vertical beam counter
	wire lineReset;
	reg [8:0] lineCounter;
	// preload data pixel counter
	reg [1:0] daCount;
	wire daCountEnable;

	always @(negedge Clk) begin
		if (colCounter == allcols) begin
			colCounter <= 9'd0; // reset columns
			HSn <= 1'b0; // start sync
			hBlank <= 1'b1; // start blank if not already running
			if (lineCounter == frameAllRows) begin
				lineCounter <= 9'd0; // reset rows
				FSn <= 1'b0; // start sync
				vBlank <= 1'b1; // start blank
			end else begin
				lineCounter <= lineCounter + 9'd1;
				if (lineCounter == 4)
					FSn <= 1'b1; // end sync
				if (lineCounter == 8)
					vBlank <= 1'b0; // end blank
			end
		end else begin
			colCounter <= colCounter + 9'd1;
			if (colCounter == leftSync)
				HSn <= 1'b1; // end sync
			if (colCounter == leftmargin)
				hBlank <= 1'b0; // end blank
			if (colCounter == rightmargin)
				hBlank <= 1'b1; // start blank
		end
		if (daCountEnable) begin
			daCount <= daCount + 2'd1;
			if (daCount == 2'b01)
				u_da0 = ~u_da0;
		end else begin
			daCount <= 2'd0;
			u_da0 = 1'b0;
		end
	end
	
	reg Clk3;
	always @(negedge Clk) begin
		Clk3 = ~Clk3;
	end

	wire alphaRowReset;
	reg [3:0] alphaRowCounter;
	always @(negedge HSn) begin
		if (alphaRowReset)
			alphaRowCounter <= 0;
		else if (activeRow)
			alphaRowCounter <= alphaRowCounter + 4'd1;
	end
	assign alphaRow = alphaRowCounter;
		
	// horizontal
	parameter leftSync = 14; // 4us duration
	parameter allcols = 227; // 64us duration (63.55)
	parameter leftmargin = 34; // 12us duration //42
	parameter rightmargin = 225; // suggested 8 cycles of front porch //225
	// vertical
	parameter activerows = 192;
	// pal
	parameter allrows = 311;// pal
	parameter topmargin = 64; //pal
	parameter toprow = 64;
	parameter bottomrow = 256; //pal
	// ntsc
	parameter allrows2 = 258;// ntsc
	parameter topmargin2 = 39; //ntsc
	parameter toprow2 = 48;
	parameter bottomrow2 = 240; //ntsc

	//parameter activecols = 128;// * 2 = 256
	parameter leftcols = 64; //
	parameter rightcols = 192; //leftcols + activecols + 1;
	parameter leftpreload = 62; //leftcols - 4;
	parameter rightpreload = 190; //rightcols - 4;

	initial begin
	   u_da0 = 1;
		colCounter = 0;
		lineCounter = 0;
		Clk3 = 0;
		alphaRowCounter = 0;
	end

	
	// vertical sync active low
	//assign FSn = ~(lineCounter[8:2] == 6'd0); 
	// 8 lines of vsync according to spec - 6847 produces nearer 40 lines...use 32 need to fix this for NTSC if I start at 16 instead of 0
	// Spectrum ULA generates just 4 lines of vsync and 8 lines of blank
	
	// horizontal sync active low
	//assign HSn = (colCounter > leftSync);

	// frame rows counter reset active high
//	assign lineReset = lineCounter == frameAllRows;
	// column counter reset active high
//	assign colReset = colCounter == allcols;
	// PAL:
	// NTSC: start lineCounter at 16?
	assign activeRow = (lineCounter > frameTopRow) && (lineCounter < frameBottomRow);
	// backporch active high
	assign BackPorch = hBlank || vBlank;
	
	assign Load = colCounter[1:0] == 0;
	assign active = activeRow && (colCounter > leftcols) && (colCounter < rightcols);
	assign daCountEnable = (activeRow && (colCounter > leftpreload));
	
	// general signals
	assign slowMode = AnG && (GMode == 3'b000);
	assign PixelClk = slowMode ? Clk3 : Clk;
	assign frameTopRow = FrameFormat ? toprow : toprow2; // FrameFormat 1=PAL/0=NTSC
	assign frameBottomRow = FrameFormat ? bottomrow : bottomrow2;
	assign frameAllRows = FrameFormat ? allrows : allrows2;
	assign alphaRowReset = alphaRowCounter == 4'b1100;
	assign DA0 = u_da0;

endmodule